`ifndef HELIX_PKG_SVH
`define HELIX_PKG_SVH

`define HELIX_INPUT_W    256
`define HELIX_CONTEXT_W  512
`define HELIX_THOUGHT_W 1024
`define HELIX_ACTION_W   256
`define HELIX_FEEDBACK_W 384

`endif // HELIX_PKG_SVH
